package sim_file_pkg;
	`include "adder_transaction.sv"
	`include "adder_generator.sv"
	`include "adder_driver.sv"
	`include "adder_monitor.sv"
	// `include "adder_coverage.sv"
	`include "scoreboard.sv"
	`include "adder_enviourment.sv"
endpackage : sim_file_pkg